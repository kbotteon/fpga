function gray_to_binary;

endfunction

function binary_to_gray;

endfunction